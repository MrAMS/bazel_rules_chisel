module dummy1;
endmodule
