module dummy0;
endmodule
